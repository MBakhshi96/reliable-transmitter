module EncryptionSBOX( Address , SBOX_out );
	input [7:0]Address;
	output [7:0]SBOX_out;

	wire [7:0]Address;
	reg [7:0]SBOX_out;
	


	always @( * )
	begin
		case ( Address )
			8'h00: SBOX_out = 8'h63;
			8'h01: SBOX_out = 8'h7c;
			8'h02: SBOX_out = 8'h77;
			8'h03: SBOX_out = 8'h7b;
			8'h04: SBOX_out = 8'hf2;
			8'h05: SBOX_out = 8'h6b;
			8'h06: SBOX_out = 8'h6f;
			8'h07: SBOX_out = 8'hc5;
			8'h08: SBOX_out = 8'h30;
			8'h09: SBOX_out = 8'h01;
			8'h0a: SBOX_out = 8'h67;
			8'h0b: SBOX_out = 8'h2b;
			8'h0c: SBOX_out = 8'hfe;
			8'h0d: SBOX_out = 8'hd7;
			8'h0e: SBOX_out = 8'hab;
			8'h0f: SBOX_out = 8'h76;
			8'h10: SBOX_out = 8'hca;
			8'h11: SBOX_out = 8'h82;
			8'h12: SBOX_out = 8'hc9;
			8'h13: SBOX_out = 8'h7d;
			8'h14: SBOX_out = 8'hfa;
			8'h15: SBOX_out = 8'h59;
			8'h16: SBOX_out = 8'h47;
			8'h17: SBOX_out = 8'hf0;
			8'h18: SBOX_out = 8'had;
			8'h19: SBOX_out = 8'hd4;
			8'h1a: SBOX_out = 8'ha2;
			8'h1b: SBOX_out = 8'haf;
			8'h1c: SBOX_out = 8'h9c;
			8'h1d: SBOX_out = 8'ha4;
			8'h1e: SBOX_out = 8'h72;
			8'h1f: SBOX_out = 8'hc0;
			8'h20: SBOX_out = 8'hb7;
			8'h21: SBOX_out = 8'hfd;
			8'h22: SBOX_out = 8'h93;
			8'h23: SBOX_out = 8'h26;
			8'h24: SBOX_out = 8'h36;
			8'h25: SBOX_out = 8'h3f;
			8'h26: SBOX_out = 8'hf7;
			8'h27: SBOX_out = 8'hcc;
			8'h28: SBOX_out = 8'h34;
			8'h29: SBOX_out = 8'ha5;
			8'h2a: SBOX_out = 8'he5;
			8'h2b: SBOX_out = 8'hf1;
			8'h2c: SBOX_out = 8'h71;
			8'h2d: SBOX_out = 8'hd8;
			8'h2e: SBOX_out = 8'h31;
			8'h2f: SBOX_out = 8'h15;
			8'h30: SBOX_out = 8'h04;
			8'h31: SBOX_out = 8'hc7;
			8'h32: SBOX_out = 8'h23;
			8'h33: SBOX_out = 8'hc3;
			8'h34: SBOX_out = 8'h18;
			8'h35: SBOX_out = 8'h96;
			8'h36: SBOX_out = 8'h05;
			8'h37: SBOX_out = 8'h9a;
			8'h38: SBOX_out = 8'h07;
			8'h39: SBOX_out = 8'h12;
			8'h3a: SBOX_out = 8'h80;
			8'h3b: SBOX_out = 8'he2;
			8'h3c: SBOX_out = 8'heb;
			8'h3d: SBOX_out = 8'h27;
			8'h3e: SBOX_out = 8'hb2;
			8'h3f: SBOX_out = 8'h75;
			8'h40: SBOX_out = 8'h09;
			8'h41: SBOX_out = 8'h83;
			8'h42: SBOX_out = 8'h2c;
			8'h43: SBOX_out = 8'h1a;
			8'h44: SBOX_out = 8'h1b;
			8'h45: SBOX_out = 8'h6e;
			8'h46: SBOX_out = 8'h5a;
			8'h47: SBOX_out = 8'ha0;
			8'h48: SBOX_out = 8'h52;
			8'h49: SBOX_out = 8'h3b;
			8'h4a: SBOX_out = 8'hd6;
			8'h4b: SBOX_out = 8'hb3;
			8'h4c: SBOX_out = 8'h29;
			8'h4d: SBOX_out = 8'he3;
			8'h4e: SBOX_out = 8'h2f;
			8'h4f: SBOX_out = 8'h84;
			8'h50: SBOX_out = 8'h53;
			8'h51: SBOX_out = 8'hd1;
			8'h52: SBOX_out = 8'h00;
			8'h53: SBOX_out = 8'hed;
			8'h54: SBOX_out = 8'h20;
			8'h55: SBOX_out = 8'hfc;
			8'h56: SBOX_out = 8'hb1;
			8'h57: SBOX_out = 8'h5b;
			8'h58: SBOX_out = 8'h6a;
			8'h59: SBOX_out = 8'hcb;
			8'h5a: SBOX_out = 8'hbe;
			8'h5b: SBOX_out = 8'h39;
			8'h5c: SBOX_out = 8'h4a;
			8'h5d: SBOX_out = 8'h4c;
			8'h5e: SBOX_out = 8'h58;
			8'h5f: SBOX_out = 8'hcf;
			8'h60: SBOX_out = 8'hd0;
			8'h61: SBOX_out = 8'hef;
			8'h62: SBOX_out = 8'haa;
			8'h63: SBOX_out = 8'hfb;
			8'h64: SBOX_out = 8'h43;
			8'h65: SBOX_out = 8'h4d;
			8'h66: SBOX_out = 8'h33;
			8'h67: SBOX_out = 8'h85;
			8'h68: SBOX_out = 8'h45;
			8'h69: SBOX_out = 8'hf9;
			8'h6a: SBOX_out = 8'h02;
			8'h6b: SBOX_out = 8'h7f;
			8'h6c: SBOX_out = 8'h50;
			8'h6d: SBOX_out = 8'h3c;
			8'h6e: SBOX_out = 8'h9f;
			8'h6f: SBOX_out = 8'ha8;
			8'h70: SBOX_out = 8'h51;
			8'h71: SBOX_out = 8'ha3;
			8'h72: SBOX_out = 8'h40;
			8'h73: SBOX_out = 8'h8f;
			8'h74: SBOX_out = 8'h92;
			8'h75: SBOX_out = 8'h9d;
			8'h76: SBOX_out = 8'h38;
			8'h77: SBOX_out = 8'hf5;
			8'h78: SBOX_out = 8'hbc;
			8'h79: SBOX_out = 8'hb6;
			8'h7a: SBOX_out = 8'hda;
			8'h7b: SBOX_out = 8'h21;
			8'h7c: SBOX_out = 8'h10;
			8'h7d: SBOX_out = 8'hff;
			8'h7e: SBOX_out = 8'hf3;
			8'h7f: SBOX_out = 8'hd2;
			8'h80: SBOX_out = 8'hcd;
			8'h81: SBOX_out = 8'h0c;
			8'h82: SBOX_out = 8'h13;
			8'h83: SBOX_out = 8'hec;
			8'h84: SBOX_out = 8'h5f;
			8'h85: SBOX_out = 8'h97;
			8'h86: SBOX_out = 8'h44;
			8'h87: SBOX_out = 8'h17;
			8'h88: SBOX_out = 8'hc4;
			8'h89: SBOX_out = 8'ha7;
			8'h8a: SBOX_out = 8'h7e;
			8'h8b: SBOX_out = 8'h3d;
			8'h8c: SBOX_out = 8'h64;
			8'h8d: SBOX_out = 8'h5d;
			8'h8e: SBOX_out = 8'h19;
			8'h8f: SBOX_out = 8'h73;
			8'h90: SBOX_out = 8'h60;
			8'h91: SBOX_out = 8'h81;
			8'h92: SBOX_out = 8'h4f;
			8'h93: SBOX_out = 8'hdc;
			8'h94: SBOX_out = 8'h22;
			8'h95: SBOX_out = 8'h2a;
			8'h96: SBOX_out = 8'h90;
			8'h97: SBOX_out = 8'h88;
			8'h98: SBOX_out = 8'h46;
			8'h99: SBOX_out = 8'hee;
			8'h9a: SBOX_out = 8'hb8;
			8'h9b: SBOX_out = 8'h14;
			8'h9c: SBOX_out = 8'hde;
			8'h9d: SBOX_out = 8'h5e;
			8'h9e: SBOX_out = 8'h0b;
			8'h9f: SBOX_out = 8'hdb;
			8'ha0: SBOX_out = 8'he0;
			8'ha1: SBOX_out = 8'h32;
			8'ha2: SBOX_out = 8'h3a;
			8'ha3: SBOX_out = 8'h0a;
			8'ha4: SBOX_out = 8'h49;
			8'ha5: SBOX_out = 8'h06;
			8'ha6: SBOX_out = 8'h24;
			8'ha7: SBOX_out = 8'h5c;
			8'ha8: SBOX_out = 8'hc2;
			8'ha9: SBOX_out = 8'hd3;
			8'haa: SBOX_out = 8'hac;
			8'hab: SBOX_out = 8'h62;
			8'hac: SBOX_out = 8'h91;
			8'had: SBOX_out = 8'h95;
			8'hae: SBOX_out = 8'he4;
			8'haf: SBOX_out = 8'h79;
			8'hb0: SBOX_out = 8'he7;
			8'hb1: SBOX_out = 8'hc8;
			8'hb2: SBOX_out = 8'h37;
			8'hb3: SBOX_out = 8'h6d;
			8'hb4: SBOX_out = 8'h8d;
			8'hb5: SBOX_out = 8'hd5;
			8'hb6: SBOX_out = 8'h4e;
			8'hb7: SBOX_out = 8'ha9;
			8'hb8: SBOX_out = 8'h6c;
			8'hb9: SBOX_out = 8'h56;
			8'hba: SBOX_out = 8'hf4;
			8'hbb: SBOX_out = 8'hea;
			8'hbc: SBOX_out = 8'h65;
			8'hbd: SBOX_out = 8'h7a;
			8'hbe: SBOX_out = 8'hae;
			8'hbf: SBOX_out = 8'h08;
			8'hc0: SBOX_out = 8'hba;
			8'hc1: SBOX_out = 8'h78;
			8'hc2: SBOX_out = 8'h25;
			8'hc3: SBOX_out = 8'h2e;
			8'hc4: SBOX_out = 8'h1c;
			8'hc5: SBOX_out = 8'ha6;
			8'hc6: SBOX_out = 8'hb4;
			8'hc7: SBOX_out = 8'hc6;
			8'hc8: SBOX_out = 8'he8;
			8'hc9: SBOX_out = 8'hdd;
			8'hca: SBOX_out = 8'h74;
			8'hcb: SBOX_out = 8'h1f;
			8'hcc: SBOX_out = 8'h4b;
			8'hcd: SBOX_out = 8'hbd;
			8'hce: SBOX_out = 8'h8b;
			8'hcf: SBOX_out = 8'h8a;
			8'hd0: SBOX_out = 8'h70;
			8'hd1: SBOX_out = 8'h3e;
			8'hd2: SBOX_out = 8'hb5;
			8'hd3: SBOX_out = 8'h66;
			8'hd4: SBOX_out = 8'h48;
			8'hd5: SBOX_out = 8'h03;
			8'hd6: SBOX_out = 8'hf6;
			8'hd7: SBOX_out = 8'h0e;
			8'hd8: SBOX_out = 8'h61;
			8'hd9: SBOX_out = 8'h35;
			8'hda: SBOX_out = 8'h57;
			8'hdb: SBOX_out = 8'hb9;
			8'hdc: SBOX_out = 8'h86;
			8'hdd: SBOX_out = 8'hc1;
			8'hde: SBOX_out = 8'h1d;
			8'hdf: SBOX_out = 8'h9e;
			8'he0: SBOX_out = 8'he1;
			8'he1: SBOX_out = 8'hf8;
			8'he2: SBOX_out = 8'h98;
			8'he3: SBOX_out = 8'h11;
			8'he4: SBOX_out = 8'h69;
			8'he5: SBOX_out = 8'hd9;
			8'he6: SBOX_out = 8'h8e;
			8'he7: SBOX_out = 8'h94;
			8'he8: SBOX_out = 8'h9b;
			8'he9: SBOX_out = 8'h1e;
			8'hea: SBOX_out = 8'h87;
			8'heb: SBOX_out = 8'he9;
			8'hec: SBOX_out = 8'hce;
			8'hed: SBOX_out = 8'h55;
			8'hee: SBOX_out = 8'h28;
			8'hef: SBOX_out = 8'hdf;
			8'hf0: SBOX_out = 8'h8c;
			8'hf1: SBOX_out = 8'ha1;
			8'hf2: SBOX_out = 8'h89;
			8'hf3: SBOX_out = 8'h0d;
			8'hf4: SBOX_out = 8'hbf;
			8'hf5: SBOX_out = 8'he6;
			8'hf6: SBOX_out = 8'h42;
			8'hf7: SBOX_out = 8'h68;
			8'hf8: SBOX_out = 8'h41;
			8'hf9: SBOX_out = 8'h99;
			8'hfa: SBOX_out = 8'h2d;
			8'hfb: SBOX_out = 8'h0f;
			8'hfc: SBOX_out = 8'hb0;
			8'hfd: SBOX_out = 8'h54;
			8'hfe: SBOX_out = 8'hbb;
			8'hff: SBOX_out = 8'h16;
		endcase
	end
	
endmodule
